module main;
	initial
		begin
			$display("DIT ME TAO");
			$finish;
		end
endmodule
