module main;
	initial
		begin
			$display("DIT ME MAY");
			$finish;
		end
endmodule